module OR_inciso2(
    output out_7,
    input out1,
    input out2,
    input out3,
    input out4,
    input out5,
    input out6
    
    
);
assign out_7 = (out1)|(out2)|(out3)|(out4)|(out5)|(out6);
endmodule

 