
module AND_inciso3(
    output out_7,
    output S_OR3,
    input Y,
    input Z,
    input K,
    input M,
    input X
);

assign noX = !X;
assign noY = !Y;
assign noZ = !Z;
assign noK = !K;
assign noM = !M;

assign out_1 = noX & noY & noM;
assign out_2 = noX & Y & K & M;
assign out_3=  noY & noZ & K;
assign out_4 = noX & noZ & K;
assign out_5 = X & noY & M;
assign out_6 = X & noZ & M;
assign S_OR3 = (out_1)|(out_2)|(out_3)|(out_4)|(out_5)|(out_6);

assign out_7 = (out_1) | (out_2) | (out_3) | (out_4) | (out_5) | (X & ~Z & M);
//assign out_7 = (~X & ~Y & ~M) | (~X & Y & K & M) | (~Y & ~Z & K) | (~X & ~Z & K) | (X & ~Y & M) | (X & ~Z & M);

endmodule     




 


