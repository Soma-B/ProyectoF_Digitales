module OR_inciso2(
    output S_OR,
    input S_1,
    input S_2,
    input S_3,
    input S_4,
    input S_5,
    input S_6,
    input S_7,
    input S_8,
    input S_9,
    input S_10,
    input S_11,
    input S_12,
    input S_13,
    input S_14    
);
assign S_OR = (S_1)|(S_2)|(S_3)|(S_4)|(S_5)|(S_6)|(S_7)|(S_7)|(S_8)|(S_9)|(S_10)|(S_11)|(S_12)|(S_13)|(S_14);
endmodule

 