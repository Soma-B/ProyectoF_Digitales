module m7(
    output out_8,
    //input noX,
    //input noY,
    //input noZ,
    //input noY,
    //input noK,
    //input noM,
   input X,
    input Y
    //input Z,
    //input K
    //input M,
    // REcordar poner noX
    
);
assign out_8 = (X)&(Y);// recordar incluir a noX
endmodule
