`include "inver.v"
`include "AND.v"
`include "OR.v"

module moduleName (
    ports
);
    
endmodule