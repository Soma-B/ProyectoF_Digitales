module f5(
    output out_7,
    input wire_out1,
    input wire_out2,
    input wire_out3,
    input wire_out4,
    input wire_out5,
    input wire_out6
    
    
);
assign out_7 = (wire_out1)|(wire_out2)|(wire_out3)|(wire_out4)|(wire_out5)|(wire_out6);// recordar incluir a noX
endmodule

 